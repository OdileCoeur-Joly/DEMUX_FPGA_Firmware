----------------------------------------------------------------------------------
-- Company       : CNRS - INSU - IRAP
-- Engineer      : Antoine CLENET / Christophe OZIOL 
-- Create Date   : 12:14:36 05/26/2015 
-- Design Name   : DRE XIFU FPGA_BOARD
-- Module Name   : Pulse_Emulator - Behavioral 
-- Project Name  : Athena XIfu DRE
-- Target Devices: Virtex 6 LX 240
-- Tool versions : ISE-14.7
-- Description: 	XXX function stored into the LUT with linear interpolation. The table must be generated using the "Function_LUT_SCRIPT.py" Python script
-- 			INSTANTIATION :
--				Size_in 	=> 22,
--				Size_out	=> 11,
-- Revision: 
-- Revision 0.1 - File Created
-- Additional Comments: 
--
---------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity LUT_func is
    Generic (
		C_Size_in			: positive;	-- 18
		C_Size_out			: positive	-- 14
		);
    Port ( 
--RESET
		RESET		: in  std_logic;
--CLOCK
		CLK			: in  std_logic;
		ENABLE_CLK	: in  std_logic;

		Func_in 	: in  unsigned(C_Size_in-1 downto 0);
		Func_out 	: out unsigned(C_Size_out-1 downto 0)
		);
end LUT_func;

--! @brief-- BLock diagrams schematics -- 
--! @detail file:work.LUT_func.Behavioral.svg
architecture Behavioral of LUT_func is

constant C_ROM_Depth 		: integer:= 11;			--  <======
constant C_Size_ROM_Sig 	: integer:= 16;		--  <======
constant C_Size_ROM_Delta	: integer:= 14;			--  <======

type LUT_func is array ((2**C_ROM_Depth)-1 downto 0) of std_logic_vector(C_Size_ROM_Sig+C_Size_ROM_Delta-1 downto 0);
constant cts_rom_data : LUT_func := (
-------------------------------------------------------------------
-- In this version of the ROM:
--   - a quarter of a period only is stored
--   - the absolute value of the Delta is stored (-1 * Delta)
--   - the sine values are stored on Size_ROM_sine bits
--   - the Delta values are stored on Size_ROM_delta bits
-------------------------------------------------------------------

0	=>	"000000000000000001010001101001",
1	=>	"000101000110100101001010000110",
2	=>	"001001101110111101000011000010",
3	=>	"001101111011001000111100101101",
4	=>	"010001101101111100110111000011",
5	=>	"010101001010000100110001111110",
6	=>	"011000010001111100101101011011",
7	=>	"011011000111101100101001010111",
8	=>	"011101101101000100100101101100",
9	=>	"100000000011111000100010011010",
10	=>	"100010001101011100011111011100",
11	=>	"100100001011001100011100110001",
12	=>	"100101111110010000011010010110",
13	=>	"100111100111101000011000001001",
14	=>	"101001001000001100010110001010",
15	=>	"101010100000110100010100010110",
16	=>	"101011110010001100010010101100",
17	=>	"101100111100111100010001001100",
18	=>	"101110000001101100001111110100",
19	=>	"101111000000111100001110100011",
20	=>	"101111111011001000001101011001",
21	=>	"110000110000101100001100010101",
22	=>	"110001100010000000001011010110",
23	=>	"110010001111011100001010011101",
24	=>	"110010111001001100001001100111",
25	=>	"110011011111101000001000110110",
26	=>	"110100000011000000001000001000",
27	=>	"110100100011100000000111011110",
28	=>	"110101000001011000000110110111",
29	=>	"110101011100110100000110010010",
30	=>	"110101110101111100000101110000",
31	=>	"110110001100111100000101010000",
32	=>	"110110100001111100000100110011",
33	=>	"110110110101001000000100010111",
34	=>	"110111000110100100000011111101",
35	=>	"110111010110011000000011100101",
36	=>	"110111100100101100000011001111",
37	=>	"110111110001101000000010111001",
38	=>	"110111111101001100000010100101",
39	=>	"111000000111100000000010010011",
40	=>	"111000010000101100000010000001",
41	=>	"111000011000110000000001110001",
42	=>	"111000011111110100000001100001",
43	=>	"111000100101111000000001010010",
44	=>	"111000101011000000000001000100",
45	=>	"111000101111010100000000110111",
46	=>	"111000110010110000000000101011",
47	=>	"111000110101011100000000011111",
48	=>	"111000110111011000000000010100",
49	=>	"111000111000101100000000001010",
50	=>	"111000111001010000000000000000",
51	=>	"111000111001010011111111110110",
52	=>	"111000111000101111111111101101",
53	=>	"111000110111100011111111100101",
54	=>	"111000110101110111111111011101",
55	=>	"111000110011101011111111010101",
56	=>	"111000110000111111111111001110",
57	=>	"111000101101110111111111000111",
58	=>	"111000101010010011111111000000",
59	=>	"111000100110010011111110111010",
60	=>	"111000100001111011111110110100",
61	=>	"111000011101001011111110101110",
62	=>	"111000011000000011111110101001",
63	=>	"111000010010100111111110100011",
64	=>	"111000001100110011111110011110",
65	=>	"111000000110101111111110011010",
66	=>	"111000000000010011111110010101",
67	=>	"110111111001100111111110010001",
68	=>	"110111110010101011111110001100",
69	=>	"110111101011011011111110001000",
70	=>	"110111100011111011111110000100",
71	=>	"110111011100001111111110000001",
72	=>	"110111010100001111111101111101",
73	=>	"110111001100000011111101111010",
74	=>	"110111000011101011111101110110",
75	=>	"110110111011000011111101110011",
76	=>	"110110110010001111111101110000",
77	=>	"110110101001001111111101101101",
78	=>	"110110100000000011111101101010",
79	=>	"110110010110101011111101100111",
80	=>	"110110001101000111111101100101",
81	=>	"110110000011011011111101100010",
82	=>	"110101111001100011111101100000",
83	=>	"110101101111011111111101011101",
84	=>	"110101100101010111111101011011",
85	=>	"110101011010111111111101011001",
86	=>	"110101010000100011111101010110",
87	=>	"110101000101111111111101010100",
88	=>	"110100111011001111111101010010",
89	=>	"110100110000010111111101010000",
90	=>	"110100100101011011111101001111",
91	=>	"110100011010010011111101001101",
92	=>	"110100001111000111111101001011",
93	=>	"110100000011110011111101001001",
94	=>	"110011111000010111111101001000",
95	=>	"110011101100110111111101000110",
96	=>	"110011100001001111111101000100",
97	=>	"110011010101011111111101000011",
98	=>	"110011001001101011111101000001",
99	=>	"110010111101101111111101000000",
100	=>	"110010110001101111111100111111",
101	=>	"110010100101101011111100111101",
102	=>	"110010011001011111111100111100",
103	=>	"110010001101001111111100111011",
104	=>	"110010000000110111111100111001",
105	=>	"110001110100011111111100111000",
106	=>	"110001100111111111111100110111",
107	=>	"110001011011011011111100110110",
108	=>	"110001001110110011111100110101",
109	=>	"110001000010000011111100110100",
110	=>	"110000110101010011111100110011",
111	=>	"110000101000011111111100110010",
112	=>	"110000011011100111111100110001",
113	=>	"110000001110100111111100110000",
114	=>	"110000000001100111111100101111",
115	=>	"101111110100100011111100101110",
116	=>	"101111100111011011111100101101",
117	=>	"101111011010001111111100101100",
118	=>	"101111001101000011111100101100",
119	=>	"101110111111101111111100101011",
120	=>	"101110110010011011111100101010",
121	=>	"101110100101000011111100101001",
122	=>	"101110010111101011111100101001",
123	=>	"101110001010001011111100101000",
124	=>	"101101111100101011111100100111",
125	=>	"101101101111000111111100100111",
126	=>	"101101100001100011111100100110",
127	=>	"101101010011111011111100100101",
128	=>	"101101000110010011111100100101",
129	=>	"101100111000100111111100100100",
130	=>	"101100101010110111111100100100",
131	=>	"101100011101000111111100100011",
132	=>	"101100001111010011111100100011",
133	=>	"101100000001011111111100100010",
134	=>	"101011110011100111111100100010",
135	=>	"101011100101101111111100100010",
136	=>	"101011010111110111111100100001",
137	=>	"101011001001111011111100100001",
138	=>	"101010111011111111111100100000",
139	=>	"101010101101111111111100100000",
140	=>	"101010100000000011111100100000",
141	=>	"101010010001111111111100011111",
142	=>	"101010000011111111111100011111",
143	=>	"101001110101111011111100011111",
144	=>	"101001100111110111111100011111",
145	=>	"101001011001110011111100011110",
146	=>	"101001001011101011111100011110",
147	=>	"101000111101100011111100011110",
148	=>	"101000101111011011111100011110",
149	=>	"101000100001010011111100011110",
150	=>	"101000010011001011111100011110",
151	=>	"101000000101000011111100011101",
152	=>	"100111110110110111111100011101",
153	=>	"100111101000101011111100011101",
154	=>	"100111011010100011111100011101",
155	=>	"100111001100010111111100011101",
156	=>	"100110111110001011111100011101",
157	=>	"100110101111111111111100011101",
158	=>	"100110100001110011111100011101",
159	=>	"100110010011100111111100011101",
160	=>	"100110000101011011111100011101",
161	=>	"100101110111001111111100011101",
162	=>	"100101101001000011111100011101",
163	=>	"100101011010111011111100011101",
164	=>	"100101001100101111111100011101",
165	=>	"100100111110100011111100011101",
166	=>	"100100110000011011111100011110",
167	=>	"100100100010001111111100011110",
168	=>	"100100010100000111111100011110",
169	=>	"100100000101111111111100011110",
170	=>	"100011110111110111111100011110",
171	=>	"100011101001101111111100011110",
172	=>	"100011011011100111111100011111",
173	=>	"100011001101100011111100011111",
174	=>	"100010111111011011111100011111",
175	=>	"100010110001010111111100011111",
176	=>	"100010100011010011111100011111",
177	=>	"100010010101010011111100100000",
178	=>	"100010000111010011111100100000",
179	=>	"100001111001010011111100100000",
180	=>	"100001101011010011111100100001",
181	=>	"100001011101010111111100100001",
182	=>	"100001001111011011111100100001",
183	=>	"100001000001011111111100100010",
184	=>	"100000110011100111111100100010",
185	=>	"100000100101101111111100100010",
186	=>	"100000010111110111111100100011",
187	=>	"100000001010000011111100100011",
188	=>	"011111111100001111111100100100",
189	=>	"011111101110011011111100100100",
190	=>	"011111100000101011111100100100",
191	=>	"011111010010111111111100100101",
192	=>	"011111000101010011111100100101",
193	=>	"011110110111100111111100100110",
194	=>	"011110101001111111111100100110",
195	=>	"011110011100010111111100100111",
196	=>	"011110001110110011111100100111",
197	=>	"011110000001001111111100101000",
198	=>	"011101110011101111111100101000",
199	=>	"011101100110001111111100101001",
200	=>	"011101011000110011111100101001",
201	=>	"011101001011011011111100101010",
202	=>	"011100111110000011111100101011",
203	=>	"011100110000101011111100101011",
204	=>	"011100100011010111111100101100",
205	=>	"011100010110000111111100101100",
206	=>	"011100001000110111111100101101",
207	=>	"011011111011101011111100101101",
208	=>	"011011101110011111111100101110",
209	=>	"011011100001011011111100101111",
210	=>	"011011010100010011111100101111",
211	=>	"011011000111010011111100110000",
212	=>	"011010111010010011111100110001",
213	=>	"011010101101010011111100110001",
214	=>	"011010100000011011111100110010",
215	=>	"011010010011100011111100110011",
216	=>	"011010000110101111111100110011",
217	=>	"011001111001111011111100110100",
218	=>	"011001101101001011111100110101",
219	=>	"011001100000011111111100110110",
220	=>	"011001010011110111111100110110",
221	=>	"011001000111001111111100110111",
222	=>	"011000111010101011111100111000",
223	=>	"011000101110001011111100111001",
224	=>	"011000100001101011111100111001",
225	=>	"011000010101010011111100111010",
226	=>	"011000001000111011111100111011",
227	=>	"010111111100100011111100111100",
228	=>	"010111110000010011111100111100",
229	=>	"010111100100000011111100111101",
230	=>	"010111010111111011111100111110",
231	=>	"010111001011110011111100111111",
232	=>	"010110111111101011111101000000",
233	=>	"010110110011101011111101000000",
234	=>	"010110100111101011111101000001",
235	=>	"010110011011110011111101000010",
236	=>	"010110001111111011111101000011",
237	=>	"010110000100000111111101000100",
238	=>	"010101111000010011111101000101",
239	=>	"010101101100100111111101000101",
240	=>	"010101100000111011111101000110",
241	=>	"010101010101010111111101000111",
242	=>	"010101001001110011111101001000",
243	=>	"010100111110010011111101001001",
244	=>	"010100110010110111111101001010",
245	=>	"010100100111011011111101001011",
246	=>	"010100011100000111111101001100",
247	=>	"010100010000110011111101001100",
248	=>	"010100000101100111111101001101",
249	=>	"010011111010011011111101001110",
250	=>	"010011101111010011111101001111",
251	=>	"010011100100001111111101010000",
252	=>	"010011011001001111111101010001",
253	=>	"010011001110010011111101010010",
254	=>	"010011000011011011111101010011",
255	=>	"010010111000100111111101010100",
256	=>	"010010101101110011111101010101",
257	=>	"010010100011000111111101010101",
258	=>	"010010011000011011111101010110",
259	=>	"010010001101110111111101010111",
260	=>	"010010000011010011111101011000",
261	=>	"010001111000110011111101011001",
262	=>	"010001101110011011111101011010",
263	=>	"010001100100000011111101011011",
264	=>	"010001011001101111111101011100",
265	=>	"010001001111011111111101011101",
266	=>	"010001000101010011111101011110",
267	=>	"010000111011001011111101011111",
268	=>	"010000110001000111111101100000",
269	=>	"010000100111000011111101100001",
270	=>	"010000011101000111111101100010",
271	=>	"010000010011001111111101100011",
272	=>	"010000001001010111111101100100",
273	=>	"001111111111100111111101100101",
274	=>	"001111110101111011111101100110",
275	=>	"001111101100001111111101100110",
276	=>	"001111100010101011111101100111",
277	=>	"001111011001000111111101101000",
278	=>	"001111001111100111111101101001",
279	=>	"001111000110001111111101101010",
280	=>	"001110111100110111111101101011",
281	=>	"001110110011100011111101101100",
282	=>	"001110101010010111111101101101",
283	=>	"001110100001001011111101101110",
284	=>	"001110011000000011111101101111",
285	=>	"001110001110111111111101110000",
286	=>	"001110000101111111111101110001",
287	=>	"001101111101000011111101110010",
288	=>	"001101110100001011111101110011",
289	=>	"001101101011010111111101110100",
290	=>	"001101100010100111111101110101",
291	=>	"001101011001111011111101110110",
292	=>	"001101010001010011111101110111",
293	=>	"001101001000101111111101111000",
294	=>	"001101000000001111111101111001",
295	=>	"001100110111110011111101111010",
296	=>	"001100101111010111111101111011",
297	=>	"001100100111000011111101111100",
298	=>	"001100011110110011111101111101",
299	=>	"001100010110100011111101111110",
300	=>	"001100001110011011111101111111",
301	=>	"001100000110010011111101111111",
302	=>	"001011111110010011111110000000",
303	=>	"001011110110010011111110000001",
304	=>	"001011101110011011111110000010",
305	=>	"001011100110100011111110000011",
306	=>	"001011011110101111111110000100",
307	=>	"001011010110111111111110000101",
308	=>	"001011001111010011111110000110",
309	=>	"001011000111101111111110000111",
310	=>	"001011000000001011111110001000",
311	=>	"001010111000100111111110001001",
312	=>	"001010110001001011111110001010",
313	=>	"001010101001110011111110001011",
314	=>	"001010100010011111111110001100",
315	=>	"001010011011001111111110001101",
316	=>	"001010010011111111111110001110",
317	=>	"001010001100110111111110001110",
318	=>	"001010000101101111111110001111",
319	=>	"001001111110101011111110010000",
320	=>	"001001110111101111111110010001",
321	=>	"001001110000110011111110010010",
322	=>	"001001101001111011111110010011",
323	=>	"001001100011000111111110010100",
324	=>	"001001011100010111111110010101",
325	=>	"001001010101101011111110010110",
326	=>	"001001001110111111111110010111",
327	=>	"001001001000011011111110010111",
328	=>	"001001000001111011111110011000",
329	=>	"001000111011011011111110011001",
330	=>	"001000110100111111111110011010",
331	=>	"001000101110100111111110011011",
332	=>	"001000101000010011111110011100",
333	=>	"001000100010000011111110011101",
334	=>	"001000011011110111111110011110",
335	=>	"001000010101101111111110011110",
336	=>	"001000001111100111111110011111",
337	=>	"001000001001100011111110100000",
338	=>	"001000000011100111111110100001",
339	=>	"000111111101101011111110100010",
340	=>	"000111110111110011111110100011",
341	=>	"000111110001111011111110100100",
342	=>	"000111101100001011111110100100",
343	=>	"000111100110011011111110100101",
344	=>	"000111100000110011111110100110",
345	=>	"000111011011001011111110100111",
346	=>	"000111010101100111111110101000",
347	=>	"000111010000000111111110101001",
348	=>	"000111001010100111111110101001",
349	=>	"000111000101001011111110101010",
350	=>	"000110111111110111111110101011",
351	=>	"000110111010100011111110101100",
352	=>	"000110110101001111111110101101",
353	=>	"000110110000000011111110101101",
354	=>	"000110101010111011111110101110",
355	=>	"000110100101110011111110101111",
356	=>	"000110100000101111111110110000",
357	=>	"000110011011101011111110110001",
358	=>	"000110010110101111111110110001",
359	=>	"000110010001110011111110110010",
360	=>	"000110001100111011111110110011",
361	=>	"000110001000000111111110110100",
362	=>	"000110000011010111111110110100",
363	=>	"000101111110100111111110110101",
364	=>	"000101111001111011111110110110",
365	=>	"000101110101010011111110110111",
366	=>	"000101110000101111111110110111",
367	=>	"000101101100001011111110111000",
368	=>	"000101100111101011111110111001",
369	=>	"000101100011001111111110111010",
370	=>	"000101011110110011111110111010",
371	=>	"000101011010011011111110111011",
372	=>	"000101010110000111111110111100",
373	=>	"000101010001110111111110111100",
374	=>	"000101001101100111111110111101",
375	=>	"000101001001011011111110111110",
376	=>	"000101000101010011111110111110",
377	=>	"000101000001001111111110111111",
378	=>	"000100111101001011111111000000",
379	=>	"000100111001001011111111000000",
380	=>	"000100110101001011111111000001",
381	=>	"000100110001001111111111000010",
382	=>	"000100101101010111111111000010",
383	=>	"000100101001011111111111000011",
384	=>	"000100100101101111111111000100",
385	=>	"000100100001111011111111000100",
386	=>	"000100011110001111111111000101",
387	=>	"000100011010100011111111000110",
388	=>	"000100010110111011111111000110",
389	=>	"000100010011010011111111000111",
390	=>	"000100001111101111111111001000",
391	=>	"000100001100001011111111001000",
392	=>	"000100001000101111111111001001",
393	=>	"000100000101001111111111001001",
394	=>	"000100000001110111111111001010",
395	=>	"000011111110011111111111001011",
396	=>	"000011111011001011111111001011",
397	=>	"000011110111110111111111001100",
398	=>	"000011110100100111111111001100",
399	=>	"000011110001010111111111001101",
400	=>	"000011101110001011111111001110",
401	=>	"000011101011000011111111001110",
402	=>	"000011100111111011111111001111",
403	=>	"000011100100110011111111001111",
404	=>	"000011100001110011111111010000",
405	=>	"000011011110101111111111010000",
406	=>	"000011011011110011111111010001",
407	=>	"000011011000110111111111010001",
408	=>	"000011010101111011111111010010",
409	=>	"000011010011000011111111010011",
410	=>	"000011010000001111111111010011",
411	=>	"000011001101011011111111010100",
412	=>	"000011001010100111111111010100",
413	=>	"000011000111111011111111010101",
414	=>	"000011000101001011111111010101",
415	=>	"000011000010011111111111010110",
416	=>	"000010111111110111111111010110",
417	=>	"000010111101001111111111010111",
418	=>	"000010111010101011111111010111",
419	=>	"000010111000000111111111011000",
420	=>	"000010110101100111111111011000",
421	=>	"000010110011000111111111011001",
422	=>	"000010110000100111111111011001",
423	=>	"000010101110001011111111011010",
424	=>	"000010101011110011111111011010",
425	=>	"000010101001011011111111011010",
426	=>	"000010100111000011111111011011",
427	=>	"000010100100101111111111011011",
428	=>	"000010100010011111111111011100",
429	=>	"000010100000001011111111011100",
430	=>	"000010011101111111111111011101",
431	=>	"000010011011101111111111011101",
432	=>	"000010011001100011111111011110",
433	=>	"000010010111011011111111011110",
434	=>	"000010010101010011111111011110",
435	=>	"000010010011001011111111011111",
436	=>	"000010010001000111111111011111",
437	=>	"000010001111000111111111100000",
438	=>	"000010001101000011111111100000",
439	=>	"000010001011000011111111100000",
440	=>	"000010001001000111111111100001",
441	=>	"000010000111001011111111100001",
442	=>	"000010000101001111111111100010",
443	=>	"000010000011010111111111100010",
444	=>	"000010000001011111111111100010",
445	=>	"000001111111100111111111100011",
446	=>	"000001111101110011111111100011",
447	=>	"000001111011111111111111100100",
448	=>	"000001111010001111111111100100",
449	=>	"000001111000011011111111100100",
450	=>	"000001110110101111111111100101",
451	=>	"000001110100111111111111100101",
452	=>	"000001110011010011111111100101",
453	=>	"000001110001101011111111100110",
454	=>	"000001101111111111111111100110",
455	=>	"000001101110010111111111100110",
456	=>	"000001101100110011111111100111",
457	=>	"000001101011001011111111100111",
458	=>	"000001101001101011111111100111",
459	=>	"000001101000000111111111101000",
460	=>	"000001100110100111111111101000",
461	=>	"000001100101000111111111101000",
462	=>	"000001100011100111111111101001",
463	=>	"000001100010001011111111101001",
464	=>	"000001100000101111111111101001",
465	=>	"000001011111010011111111101010",
466	=>	"000001011101110111111111101010",
467	=>	"000001011100011111111111101010",
468	=>	"000001011011000111111111101010",
469	=>	"000001011001110011111111101011",
470	=>	"000001011000011111111111101011",
471	=>	"000001010111001011111111101011",
472	=>	"000001010101110111111111101100",
473	=>	"000001010100100111111111101100",
474	=>	"000001010011010011111111101100",
475	=>	"000001010010000111111111101100",
476	=>	"000001010000110111111111101101",
477	=>	"000001001111101011111111101101",
478	=>	"000001001110011111111111101101",
479	=>	"000001001101010011111111101101",
480	=>	"000001001100000111111111101110",
481	=>	"000001001010111111111111101110",
482	=>	"000001001001110111111111101110",
483	=>	"000001001000101111111111101110",
484	=>	"000001000111101011111111101111",
485	=>	"000001000110100011111111101111",
486	=>	"000001000101011111111111101111",
487	=>	"000001000100011111111111101111",
488	=>	"000001000011011011111111110000",
489	=>	"000001000010011011111111110000",
490	=>	"000001000001010111111111110000",
491	=>	"000001000000011011111111110000",
492	=>	"000000111111011011111111110001",
493	=>	"000000111110011011111111110001",
494	=>	"000000111101011111111111110001",
495	=>	"000000111100100011111111110001",
496	=>	"000000111011100111111111110001",
497	=>	"000000111010101111111111110010",
498	=>	"000000111001110011111111110010",
499	=>	"000000111000111011111111110010",
500	=>	"000000111000000011111111110010",
501	=>	"000000110111001111111111110010",
502	=>	"000000110110010111111111110011",
503	=>	"000000110101100011111111110011",
504	=>	"000000110100101011111111110011",
505	=>	"000000110011110111111111110011",
506	=>	"000000110011000111111111110011",
507	=>	"000000110010010011111111110100",
508	=>	"000000110001011111111111110100",
509	=>	"000000110000101111111111110100",
510	=>	"000000101111111111111111110100",
511	=>	"000000101111001111111111110100",
512	=>	"000000101110011111111111110100",
513	=>	"000000101101110011111111110101",
514	=>	"000000101101000011111111110101",
515	=>	"000000101100010111111111110101",
516	=>	"000000101011101011111111110101",
517	=>	"000000101010111111111111110101",
518	=>	"000000101010010011111111110101",
519	=>	"000000101001101011111111110110",
520	=>	"000000101000111111111111110110",
521	=>	"000000101000010111111111110110",
522	=>	"000000100111101111111111110110",
523	=>	"000000100111000111111111110110",
524	=>	"000000100110011111111111110110",
525	=>	"000000100101110111111111110110",
526	=>	"000000100101010011111111110111",
527	=>	"000000100100101111111111110111",
528	=>	"000000100100000111111111110111",
529	=>	"000000100011100011111111110111",
530	=>	"000000100010111111111111110111",
531	=>	"000000100010011011111111110111",
532	=>	"000000100001111011111111110111",
533	=>	"000000100001010111111111111000",
534	=>	"000000100000110011111111111000",
535	=>	"000000100000010011111111111000",
536	=>	"000000011111110011111111111000",
537	=>	"000000011111010011111111111000",
538	=>	"000000011110110011111111111000",
539	=>	"000000011110010011111111111000",
540	=>	"000000011101110011111111111000",
541	=>	"000000011101010111111111111000",
542	=>	"000000011100110111111111111001",
543	=>	"000000011100011011111111111001",
544	=>	"000000011011111011111111111001",
545	=>	"000000011011011111111111111001",
546	=>	"000000011011000011111111111001",
547	=>	"000000011010100111111111111001",
548	=>	"000000011010001011111111111001",
549	=>	"000000011001110011111111111001",
550	=>	"000000011001010111111111111001",
551	=>	"000000011000111111111111111010",
552	=>	"000000011000100011111111111010",
553	=>	"000000011000001011111111111010",
554	=>	"000000010111110011111111111010",
555	=>	"000000010111010111111111111010",
556	=>	"000000010110111111111111111010",
557	=>	"000000010110100111111111111010",
558	=>	"000000010110010011111111111010",
559	=>	"000000010101111011111111111010",
560	=>	"000000010101100011111111111010",
561	=>	"000000010101001111111111111010",
562	=>	"000000010100110111111111111011",
563	=>	"000000010100100011111111111011",
564	=>	"000000010100001011111111111011",
565	=>	"000000010011110111111111111011",
566	=>	"000000010011100011111111111011",
567	=>	"000000010011001111111111111011",
568	=>	"000000010010111011111111111011",
569	=>	"000000010010100111111111111011",
570	=>	"000000010010010011111111111011",
571	=>	"000000010001111111111111111011",
572	=>	"000000010001101011111111111011",
573	=>	"000000010001011011111111111011",
574	=>	"000000010001000111111111111100",
575	=>	"000000010000110111111111111100",
576	=>	"000000010000100011111111111100",
577	=>	"000000010000010011111111111100",
578	=>	"000000010000000011111111111100",
579	=>	"000000001111101111111111111100",
580	=>	"000000001111011111111111111100",
581	=>	"000000001111001111111111111100",
582	=>	"000000001110111111111111111100",
583	=>	"000000001110101111111111111100",
584	=>	"000000001110011111111111111100",
585	=>	"000000001110010011111111111100",
586	=>	"000000001110000011111111111100",
587	=>	"000000001101110011111111111100",
588	=>	"000000001101100011111111111100",
589	=>	"000000001101010111111111111100",
590	=>	"000000001101000111111111111101",
591	=>	"000000001100111011111111111101",
592	=>	"000000001100101011111111111101",
593	=>	"000000001100011111111111111101",
594	=>	"000000001100010011111111111101",
595	=>	"000000001100000011111111111101",
596	=>	"000000001011110111111111111101",
597	=>	"000000001011101011111111111101",
598	=>	"000000001011011111111111111101",
599	=>	"000000001011010011111111111101",
600	=>	"000000001011000111111111111101",
601	=>	"000000001010111011111111111101",
602	=>	"000000001010101111111111111101",
603	=>	"000000001010100011111111111101",
604	=>	"000000001010010111111111111101",
605	=>	"000000001010001111111111111101",
606	=>	"000000001010000011111111111101",
607	=>	"000000001001110111111111111101",
608	=>	"000000001001101111111111111101",
609	=>	"000000001001100011111111111101",
610	=>	"000000001001010111111111111101",
611	=>	"000000001001001111111111111110",
612	=>	"000000001001000011111111111110",
613	=>	"000000001000111011111111111110",
614	=>	"000000001000110011111111111110",
615	=>	"000000001000100111111111111110",
616	=>	"000000001000011111111111111110",
617	=>	"000000001000010111111111111110",
618	=>	"000000001000001011111111111110",
619	=>	"000000001000000011111111111110",
620	=>	"000000000111111011111111111110",
621	=>	"000000000111110011111111111110",
622	=>	"000000000111101011111111111110",
623	=>	"000000000111100011111111111110",
624	=>	"000000000111011011111111111110",
625	=>	"000000000111010011111111111110",
626	=>	"000000000111001011111111111110",
627	=>	"000000000111000011111111111110",
628	=>	"000000000110111011111111111110",
629	=>	"000000000110110011111111111110",
630	=>	"000000000110101011111111111110",
631	=>	"000000000110100011111111111110",
632	=>	"000000000110011111111111111110",
633	=>	"000000000110010111111111111110",
634	=>	"000000000110001111111111111110",
635	=>	"000000000110001011111111111110",
636	=>	"000000000110000011111111111110",
637	=>	"000000000101111011111111111110",
638	=>	"000000000101110111111111111110",
639	=>	"000000000101101111111111111110",
640	=>	"000000000101100111111111111110",
641	=>	"000000000101100011111111111110",
642	=>	"000000000101011011111111111111",
643	=>	"000000000101010111111111111111",
644	=>	"000000000101010011111111111111",
645	=>	"000000000101001011111111111111",
646	=>	"000000000101000111111111111111",
647	=>	"000000000100111111111111111111",
648	=>	"000000000100111011111111111111",
649	=>	"000000000100110111111111111111",
650	=>	"000000000100101111111111111111",
651	=>	"000000000100101011111111111111",
652	=>	"000000000100100111111111111111",
653	=>	"000000000100011111111111111111",
654	=>	"000000000100011011111111111111",
655	=>	"000000000100010111111111111111",
656	=>	"000000000100010011111111111111",
657	=>	"000000000100001111111111111111",
658	=>	"000000000100001011111111111111",
659	=>	"000000000100000011111111111111",
660	=>	"000000000011111111111111111111",
661	=>	"000000000011111011111111111111",
662	=>	"000000000011110111111111111111",
663	=>	"000000000011110011111111111111",
664	=>	"000000000011101111111111111111",
665	=>	"000000000011101011111111111111",
666	=>	"000000000011100111111111111111",
667	=>	"000000000011100011111111111111",
668	=>	"000000000011011111111111111111",
669	=>	"000000000011011011111111111111",
670	=>	"000000000011010111111111111111",
671	=>	"000000000011010011111111111111",
672	=>	"000000000011001111111111111111",
673	=>	"000000000011001011111111111111",
674	=>	"000000000011001011111111111111",
675	=>	"000000000011000111111111111111",
676	=>	"000000000011000011111111111111",
677	=>	"000000000010111111111111111111",
678	=>	"000000000010111011111111111111",
679	=>	"000000000010110111111111111111",
680	=>	"000000000010110111111111111111",
681	=>	"000000000010110011111111111111",
682	=>	"000000000010101111111111111111",
683	=>	"000000000010101011111111111111",
684	=>	"000000000010101011111111111111",
685	=>	"000000000010100111111111111111",
686	=>	"000000000010100011111111111111",
687	=>	"000000000010011111111111111111",
688	=>	"000000000010011111111111111111",
689	=>	"000000000010011011111111111111",
690	=>	"000000000010010111111111111111",
691	=>	"000000000010010111111111111111",
692	=>	"000000000010010011111111111111",
693	=>	"000000000010010011111111111111",
694	=>	"000000000010001111111111111111",
695	=>	"000000000010001011111111111111",
696	=>	"000000000010001011111111111111",
697	=>	"000000000010000111111111111111",
698	=>	"000000000010000111111111111111",
699	=>	"000000000010000011111111111111",
700	=>	"000000000001111111111111111111",
701	=>	"000000000001111111111111111111",
702	=>	"000000000001111011111111111111",
703	=>	"000000000001111011111111111111",
704	=>	"000000000001110111111111111111",
705	=>	"000000000001110111111111111111",
706	=>	"000000000001110000000000000000",
707	=>	"000000000001110000000000000000",
708	=>	"000000000001101100000000000000",
709	=>	"000000000001101100000000000000",
710	=>	"000000000001101000000000000000",
711	=>	"000000000001101000000000000000",
712	=>	"000000000001100100000000000000",
713	=>	"000000000001100100000000000000",
714	=>	"000000000001100000000000000000",
715	=>	"000000000001100000000000000000",
716	=>	"000000000001100000000000000000",
717	=>	"000000000001011100000000000000",
718	=>	"000000000001011100000000000000",
719	=>	"000000000001011000000000000000",
720	=>	"000000000001011000000000000000",
721	=>	"000000000001011000000000000000",
722	=>	"000000000001010100000000000000",
723	=>	"000000000001010100000000000000",
724	=>	"000000000001010000000000000000",
725	=>	"000000000001010000000000000000",
726	=>	"000000000001010000000000000000",
727	=>	"000000000001001100000000000000",
728	=>	"000000000001001100000000000000",
729	=>	"000000000001001100000000000000",
730	=>	"000000000001001000000000000000",
731	=>	"000000000001001000000000000000",
732	=>	"000000000001001000000000000000",
733	=>	"000000000001000100000000000000",
734	=>	"000000000001000100000000000000",
735	=>	"000000000001000100000000000000",
736	=>	"000000000001000100000000000000",
737	=>	"000000000001000000000000000000",
738	=>	"000000000001000000000000000000",
739	=>	"000000000001000000000000000000",
740	=>	"000000000000111100000000000000",
741	=>	"000000000000111100000000000000",
742	=>	"000000000000111100000000000000",
743	=>	"000000000000111100000000000000",
744	=>	"000000000000111000000000000000",
745	=>	"000000000000111000000000000000",
746	=>	"000000000000111000000000000000",
747	=>	"000000000000111000000000000000",
748	=>	"000000000000110100000000000000",
749	=>	"000000000000110100000000000000",
750	=>	"000000000000110100000000000000",
751	=>	"000000000000110100000000000000",
752	=>	"000000000000110000000000000000",
753	=>	"000000000000110000000000000000",
754	=>	"000000000000110000000000000000",
755	=>	"000000000000110000000000000000",
756	=>	"000000000000110000000000000000",
757	=>	"000000000000101100000000000000",
758	=>	"000000000000101100000000000000",
759	=>	"000000000000101100000000000000",
760	=>	"000000000000101100000000000000",
761	=>	"000000000000101100000000000000",
762	=>	"000000000000101000000000000000",
763	=>	"000000000000101000000000000000",
764	=>	"000000000000101000000000000000",
765	=>	"000000000000101000000000000000",
766	=>	"000000000000101000000000000000",
767	=>	"000000000000100100000000000000",
768	=>	"000000000000100100000000000000",
769	=>	"000000000000100100000000000000",
770	=>	"000000000000100100000000000000",
771	=>	"000000000000100100000000000000",
772	=>	"000000000000100100000000000000",
773	=>	"000000000000100100000000000000",
774	=>	"000000000000100000000000000000",
775	=>	"000000000000100000000000000000",
776	=>	"000000000000100000000000000000",
777	=>	"000000000000100000000000000000",
778	=>	"000000000000100000000000000000",
779	=>	"000000000000100000000000000000",
780	=>	"000000000000011100000000000000",
781	=>	"000000000000011100000000000000",
782	=>	"000000000000011100000000000000",
783	=>	"000000000000011100000000000000",
784	=>	"000000000000011100000000000000",
785	=>	"000000000000011100000000000000",
786	=>	"000000000000011100000000000000",
787	=>	"000000000000011100000000000000",
788	=>	"000000000000011000000000000000",
789	=>	"000000000000011000000000000000",
790	=>	"000000000000011000000000000000",
791	=>	"000000000000011000000000000000",
792	=>	"000000000000011000000000000000",
793	=>	"000000000000011000000000000000",
794	=>	"000000000000011000000000000000",
795	=>	"000000000000011000000000000000",
796	=>	"000000000000011000000000000000",
797	=>	"000000000000011000000000000000",
798	=>	"000000000000010100000000000000",
799	=>	"000000000000010100000000000000",
800	=>	"000000000000010100000000000000",
801	=>	"000000000000010100000000000000",
802	=>	"000000000000010100000000000000",
803	=>	"000000000000010100000000000000",
804	=>	"000000000000010100000000000000",
805	=>	"000000000000010100000000000000",
806	=>	"000000000000010100000000000000",
807	=>	"000000000000010100000000000000",
808	=>	"000000000000010100000000000000",
809	=>	"000000000000010000000000000000",
810	=>	"000000000000010000000000000000",
811	=>	"000000000000010000000000000000",
812	=>	"000000000000010000000000000000",
813	=>	"000000000000010000000000000000",
814	=>	"000000000000010000000000000000",
815	=>	"000000000000010000000000000000",
816	=>	"000000000000010000000000000000",
817	=>	"000000000000010000000000000000",
818	=>	"000000000000010000000000000000",
819	=>	"000000000000010000000000000000",
820	=>	"000000000000010000000000000000",
821	=>	"000000000000010000000000000000",
822	=>	"000000000000001100000000000000",
823	=>	"000000000000001100000000000000",
824	=>	"000000000000001100000000000000",
825	=>	"000000000000001100000000000000",
826	=>	"000000000000001100000000000000",
827	=>	"000000000000001100000000000000",
828	=>	"000000000000001100000000000000",
829	=>	"000000000000001100000000000000",
830	=>	"000000000000001100000000000000",
831	=>	"000000000000001100000000000000",
832	=>	"000000000000001100000000000000",
833	=>	"000000000000001100000000000000",
834	=>	"000000000000001100000000000000",
835	=>	"000000000000001100000000000000",
836	=>	"000000000000001100000000000000",
837	=>	"000000000000001100000000000000",
838	=>	"000000000000001100000000000000",
839	=>	"000000000000001100000000000000",
840	=>	"000000000000001100000000000000",
841	=>	"000000000000001000000000000000",
842	=>	"000000000000001000000000000000",
843	=>	"000000000000001000000000000000",
844	=>	"000000000000001000000000000000",
845	=>	"000000000000001000000000000000",
846	=>	"000000000000001000000000000000",
847	=>	"000000000000001000000000000000",
848	=>	"000000000000001000000000000000",
849	=>	"000000000000001000000000000000",
850	=>	"000000000000001000000000000000",
851	=>	"000000000000001000000000000000",
852	=>	"000000000000001000000000000000",
853	=>	"000000000000001000000000000000",
854	=>	"000000000000001000000000000000",
855	=>	"000000000000001000000000000000",
856	=>	"000000000000001000000000000000",
857	=>	"000000000000001000000000000000",
858	=>	"000000000000001000000000000000",
859	=>	"000000000000001000000000000000",
860	=>	"000000000000001000000000000000",
861	=>	"000000000000001000000000000000",
862	=>	"000000000000001000000000000000",
863	=>	"000000000000001000000000000000",
864	=>	"000000000000001000000000000000",
865	=>	"000000000000001000000000000000",
866	=>	"000000000000001000000000000000",
867	=>	"000000000000001000000000000000",
868	=>	"000000000000000100000000000000",
869	=>	"000000000000000100000000000000",
870	=>	"000000000000000100000000000000",
871	=>	"000000000000000100000000000000",
872	=>	"000000000000000100000000000000",
873	=>	"000000000000000100000000000000",
874	=>	"000000000000000100000000000000",
875	=>	"000000000000000100000000000000",
876	=>	"000000000000000100000000000000",
877	=>	"000000000000000100000000000000",
878	=>	"000000000000000100000000000000",
879	=>	"000000000000000100000000000000",
880	=>	"000000000000000100000000000000",
881	=>	"000000000000000100000000000000",
882	=>	"000000000000000100000000000000",
883	=>	"000000000000000100000000000000",
884	=>	"000000000000000100000000000000",
885	=>	"000000000000000100000000000000",
886	=>	"000000000000000100000000000000",
887	=>	"000000000000000100000000000000",
888	=>	"000000000000000100000000000000",
889	=>	"000000000000000100000000000000",
890	=>	"000000000000000100000000000000",
891	=>	"000000000000000100000000000000",
892	=>	"000000000000000100000000000000",
893	=>	"000000000000000100000000000000",
894	=>	"000000000000000100000000000000",
895	=>	"000000000000000100000000000000",
896	=>	"000000000000000100000000000000",
897	=>	"000000000000000100000000000000",
898	=>	"000000000000000100000000000000",
899	=>	"000000000000000100000000000000",
900	=>	"000000000000000100000000000000",
901	=>	"000000000000000100000000000000",
902	=>	"000000000000000100000000000000",
903	=>	"000000000000000100000000000000",
904	=>	"000000000000000100000000000000",
905	=>	"000000000000000100000000000000",
906	=>	"000000000000000100000000000000",
907	=>	"000000000000000100000000000000",
908	=>	"000000000000000100000000000000",
909	=>	"000000000000000100000000000000",
910	=>	"000000000000000100000000000000",
911	=>	"000000000000000100000000000000",
912	=>	"000000000000000100000000000000",
913	=>	"000000000000000100000000000000",
914	=>	"000000000000000100000000000000",
915	=>	"000000000000000100000000000000",
916	=>	"000000000000000100000000000000",
917	=>	"000000000000000100000000000000",
918	=>	"000000000000000100000000000000",
919	=>	"000000000000000100000000000000",
920	=>	"000000000000000100000000000000",
921	=>	"000000000000000100000000000000",
922	=>	"000000000000000100000000000000",
923	=>	"000000000000000100000000000000",
924	=>	"000000000000000100000000000000",
925	=>	"000000000000000100000000000000",
926	=>	"000000000000000100000000000000",
927	=>	"000000000000000100000000000000",
928	=>	"000000000000000000000000000000",
929	=>	"000000000000000000000000000000",
930	=>	"000000000000000000000000000000",
931	=>	"000000000000000000000000000000",
932	=>	"000000000000000000000000000000",
933	=>	"000000000000000000000000000000",
934	=>	"000000000000000000000000000000",
935	=>	"000000000000000000000000000000",
936	=>	"000000000000000000000000000000",
937	=>	"000000000000000000000000000000",
938	=>	"000000000000000000000000000000",
939	=>	"000000000000000000000000000000",
940	=>	"000000000000000000000000000000",
941	=>	"000000000000000000000000000000",
942	=>	"000000000000000000000000000000",
943	=>	"000000000000000000000000000000",
944	=>	"000000000000000000000000000000",
945	=>	"000000000000000000000000000000",
946	=>	"000000000000000000000000000000",
947	=>	"000000000000000000000000000000",
948	=>	"000000000000000000000000000000",
949	=>	"000000000000000000000000000000",
950	=>	"000000000000000000000000000000",
951	=>	"000000000000000000000000000000",
952	=>	"000000000000000000000000000000",
953	=>	"000000000000000000000000000000",
954	=>	"000000000000000000000000000000",
955	=>	"000000000000000000000000000000",
956	=>	"000000000000000000000000000000",
957	=>	"000000000000000000000000000000",
958	=>	"000000000000000000000000000000",
959	=>	"000000000000000000000000000000",
960	=>	"000000000000000000000000000000",
961	=>	"000000000000000000000000000000",
962	=>	"000000000000000000000000000000",
963	=>	"000000000000000000000000000000",
964	=>	"000000000000000000000000000000",
965	=>	"000000000000000000000000000000",
966	=>	"000000000000000000000000000000",
967	=>	"000000000000000000000000000000",
968	=>	"000000000000000000000000000000",
969	=>	"000000000000000000000000000000",
970	=>	"000000000000000000000000000000",
971	=>	"000000000000000000000000000000",
972	=>	"000000000000000000000000000000",
973	=>	"000000000000000000000000000000",
974	=>	"000000000000000000000000000000",
975	=>	"000000000000000000000000000000",
976	=>	"000000000000000000000000000000",
977	=>	"000000000000000000000000000000",
978	=>	"000000000000000000000000000000",
979	=>	"000000000000000000000000000000",
980	=>	"000000000000000000000000000000",
981	=>	"000000000000000000000000000000",
982	=>	"000000000000000000000000000000",
983	=>	"000000000000000000000000000000",
984	=>	"000000000000000000000000000000",
985	=>	"000000000000000000000000000000",
986	=>	"000000000000000000000000000000",
987	=>	"000000000000000000000000000000",
988	=>	"000000000000000000000000000000",
989	=>	"000000000000000000000000000000",
990	=>	"000000000000000000000000000000",
991	=>	"000000000000000000000000000000",
992	=>	"000000000000000000000000000000",
993	=>	"000000000000000000000000000000",
994	=>	"000000000000000000000000000000",
995	=>	"000000000000000000000000000000",
996	=>	"000000000000000000000000000000",
997	=>	"000000000000000000000000000000",
998	=>	"000000000000000000000000000000",
999	=>	"000000000000000000000000000000",
1000	=>	"000000000000000000000000000000",
1001	=>	"000000000000000000000000000000",
1002	=>	"000000000000000000000000000000",
1003	=>	"000000000000000000000000000000",
1004	=>	"000000000000000000000000000000",
1005	=>	"000000000000000000000000000000",
1006	=>	"000000000000000000000000000000",
1007	=>	"000000000000000000000000000000",
1008	=>	"000000000000000000000000000000",
1009	=>	"000000000000000000000000000000",
1010	=>	"000000000000000000000000000000",
1011	=>	"000000000000000000000000000000",
1012	=>	"000000000000000000000000000000",
1013	=>	"000000000000000000000000000000",
1014	=>	"000000000000000000000000000000",
1015	=>	"000000000000000000000000000000",
1016	=>	"000000000000000000000000000000",
1017	=>	"000000000000000000000000000000",
1018	=>	"000000000000000000000000000000",
1019	=>	"000000000000000000000000000000",
1020	=>	"000000000000000000000000000000",
1021	=>	"000000000000000000000000000000",
1022	=>	"000000000000000000000000000000",
1023	=>	"000000000000000000000000000000",
1024	=>	"000000000000000000000000000000",
1025	=>	"000000000000000000000000000000",
1026	=>	"000000000000000000000000000000",
1027	=>	"000000000000000000000000000000",
1028	=>	"000000000000000000000000000000",
1029	=>	"000000000000000000000000000000",
1030	=>	"000000000000000000000000000000",
1031	=>	"000000000000000000000000000000",
1032	=>	"000000000000000000000000000000",
1033	=>	"000000000000000000000000000000",
1034	=>	"000000000000000000000000000000",
1035	=>	"000000000000000000000000000000",
1036	=>	"000000000000000000000000000000",
1037	=>	"000000000000000000000000000000",
1038	=>	"000000000000000000000000000000",
1039	=>	"000000000000000000000000000000",
1040	=>	"000000000000000000000000000000",
1041	=>	"000000000000000000000000000000",
1042	=>	"000000000000000000000000000000",
1043	=>	"000000000000000000000000000000",
1044	=>	"000000000000000000000000000000",
1045	=>	"000000000000000000000000000000",
1046	=>	"000000000000000000000000000000",
1047	=>	"000000000000000000000000000000",
1048	=>	"000000000000000000000000000000",
1049	=>	"000000000000000000000000000000",
1050	=>	"000000000000000000000000000000",
1051	=>	"000000000000000000000000000000",
1052	=>	"000000000000000000000000000000",
1053	=>	"000000000000000000000000000000",
1054	=>	"000000000000000000000000000000",
1055	=>	"000000000000000000000000000000",
1056	=>	"000000000000000000000000000000",
1057	=>	"000000000000000000000000000000",
1058	=>	"000000000000000000000000000000",
1059	=>	"000000000000000000000000000000",
1060	=>	"000000000000000000000000000000",
1061	=>	"000000000000000000000000000000",
1062	=>	"000000000000000000000000000000",
1063	=>	"000000000000000000000000000000",
1064	=>	"000000000000000000000000000000",
1065	=>	"000000000000000000000000000000",
1066	=>	"000000000000000000000000000000",
1067	=>	"000000000000000000000000000000",
1068	=>	"000000000000000000000000000000",
1069	=>	"000000000000000000000000000000",
1070	=>	"000000000000000000000000000000",
1071	=>	"000000000000000000000000000000",
1072	=>	"000000000000000000000000000000",
1073	=>	"000000000000000000000000000000",
1074	=>	"000000000000000000000000000000",
1075	=>	"000000000000000000000000000000",
1076	=>	"000000000000000000000000000000",
1077	=>	"000000000000000000000000000000",
1078	=>	"000000000000000000000000000000",
1079	=>	"000000000000000000000000000000",
1080	=>	"000000000000000000000000000000",
1081	=>	"000000000000000000000000000000",
1082	=>	"000000000000000000000000000000",
1083	=>	"000000000000000000000000000000",
1084	=>	"000000000000000000000000000000",
1085	=>	"000000000000000000000000000000",
1086	=>	"000000000000000000000000000000",
1087	=>	"000000000000000000000000000000",
1088	=>	"000000000000000000000000000000",
1089	=>	"000000000000000000000000000000",
1090	=>	"000000000000000000000000000000",
1091	=>	"000000000000000000000000000000",
1092	=>	"000000000000000000000000000000",
1093	=>	"000000000000000000000000000000",
1094	=>	"000000000000000000000000000000",
1095	=>	"000000000000000000000000000000",
1096	=>	"000000000000000000000000000000",
1097	=>	"000000000000000000000000000000",
1098	=>	"000000000000000000000000000000",
1099	=>	"000000000000000000000000000000",
1100	=>	"000000000000000000000000000000",
1101	=>	"000000000000000000000000000000",
1102	=>	"000000000000000000000000000000",
1103	=>	"000000000000000000000000000000",
1104	=>	"000000000000000000000000000000",
1105	=>	"000000000000000000000000000000",
1106	=>	"000000000000000000000000000000",
1107	=>	"000000000000000000000000000000",
1108	=>	"000000000000000000000000000000",
1109	=>	"000000000000000000000000000000",
1110	=>	"000000000000000000000000000000",
1111	=>	"000000000000000000000000000000",
1112	=>	"000000000000000000000000000000",
1113	=>	"000000000000000000000000000000",
1114	=>	"000000000000000000000000000000",
1115	=>	"000000000000000000000000000000",
1116	=>	"000000000000000000000000000000",
1117	=>	"000000000000000000000000000000",
1118	=>	"000000000000000000000000000000",
1119	=>	"000000000000000000000000000000",
1120	=>	"000000000000000000000000000000",
1121	=>	"000000000000000000000000000000",
1122	=>	"000000000000000000000000000000",
1123	=>	"000000000000000000000000000000",
1124	=>	"000000000000000000000000000000",
1125	=>	"000000000000000000000000000000",
1126	=>	"000000000000000000000000000000",
1127	=>	"000000000000000000000000000000",
1128	=>	"000000000000000000000000000000",
1129	=>	"000000000000000000000000000000",
1130	=>	"000000000000000000000000000000",
1131	=>	"000000000000000000000000000000",
1132	=>	"000000000000000000000000000000",
1133	=>	"000000000000000000000000000000",
1134	=>	"000000000000000000000000000000",
1135	=>	"000000000000000000000000000000",
1136	=>	"000000000000000000000000000000",
1137	=>	"000000000000000000000000000000",
1138	=>	"000000000000000000000000000000",
1139	=>	"000000000000000000000000000000",
1140	=>	"000000000000000000000000000000",
1141	=>	"000000000000000000000000000000",
1142	=>	"000000000000000000000000000000",
1143	=>	"000000000000000000000000000000",
1144	=>	"000000000000000000000000000000",
1145	=>	"000000000000000000000000000000",
1146	=>	"000000000000000000000000000000",
1147	=>	"000000000000000000000000000000",
1148	=>	"000000000000000000000000000000",
1149	=>	"000000000000000000000000000000",
1150	=>	"000000000000000000000000000000",
1151	=>	"000000000000000000000000000000",
1152	=>	"000000000000000000000000000000",
1153	=>	"000000000000000000000000000000",
1154	=>	"000000000000000000000000000000",
1155	=>	"000000000000000000000000000000",
1156	=>	"000000000000000000000000000000",
1157	=>	"000000000000000000000000000000",
1158	=>	"000000000000000000000000000000",
1159	=>	"000000000000000000000000000000",
1160	=>	"000000000000000000000000000000",
1161	=>	"000000000000000000000000000000",
1162	=>	"000000000000000000000000000000",
1163	=>	"000000000000000000000000000000",
1164	=>	"000000000000000000000000000000",
1165	=>	"000000000000000000000000000000",
1166	=>	"000000000000000000000000000000",
1167	=>	"000000000000000000000000000000",
1168	=>	"000000000000000000000000000000",
1169	=>	"000000000000000000000000000000",
1170	=>	"000000000000000000000000000000",
1171	=>	"000000000000000000000000000000",
1172	=>	"000000000000000000000000000000",
1173	=>	"000000000000000000000000000000",
1174	=>	"000000000000000000000000000000",
1175	=>	"000000000000000000000000000000",
1176	=>	"000000000000000000000000000000",
1177	=>	"000000000000000000000000000000",
1178	=>	"000000000000000000000000000000",
1179	=>	"000000000000000000000000000000",
1180	=>	"000000000000000000000000000000",
1181	=>	"000000000000000000000000000000",
1182	=>	"000000000000000000000000000000",
1183	=>	"000000000000000000000000000000",
1184	=>	"000000000000000000000000000000",
1185	=>	"000000000000000000000000000000",
1186	=>	"000000000000000000000000000000",
1187	=>	"000000000000000000000000000000",
1188	=>	"000000000000000000000000000000",
1189	=>	"000000000000000000000000000000",
1190	=>	"000000000000000000000000000000",
1191	=>	"000000000000000000000000000000",
1192	=>	"000000000000000000000000000000",
1193	=>	"000000000000000000000000000000",
1194	=>	"000000000000000000000000000000",
1195	=>	"000000000000000000000000000000",
1196	=>	"000000000000000000000000000000",
1197	=>	"000000000000000000000000000000",
1198	=>	"000000000000000000000000000000",
1199	=>	"000000000000000000000000000000",
1200	=>	"000000000000000000000000000000",
1201	=>	"000000000000000000000000000000",
1202	=>	"000000000000000000000000000000",
1203	=>	"000000000000000000000000000000",
1204	=>	"000000000000000000000000000000",
1205	=>	"000000000000000000000000000000",
1206	=>	"000000000000000000000000000000",
1207	=>	"000000000000000000000000000000",
1208	=>	"000000000000000000000000000000",
1209	=>	"000000000000000000000000000000",
1210	=>	"000000000000000000000000000000",
1211	=>	"000000000000000000000000000000",
1212	=>	"000000000000000000000000000000",
1213	=>	"000000000000000000000000000000",
1214	=>	"000000000000000000000000000000",
1215	=>	"000000000000000000000000000000",
1216	=>	"000000000000000000000000000000",
1217	=>	"000000000000000000000000000000",
1218	=>	"000000000000000000000000000000",
1219	=>	"000000000000000000000000000000",
1220	=>	"000000000000000000000000000000",
1221	=>	"000000000000000000000000000000",
1222	=>	"000000000000000000000000000000",
1223	=>	"000000000000000000000000000000",
1224	=>	"000000000000000000000000000000",
1225	=>	"000000000000000000000000000000",
1226	=>	"000000000000000000000000000000",
1227	=>	"000000000000000000000000000000",
1228	=>	"000000000000000000000000000000",
1229	=>	"000000000000000000000000000000",
1230	=>	"000000000000000000000000000000",
1231	=>	"000000000000000000000000000000",
1232	=>	"000000000000000000000000000000",
1233	=>	"000000000000000000000000000000",
1234	=>	"000000000000000000000000000000",
1235	=>	"000000000000000000000000000000",
1236	=>	"000000000000000000000000000000",
1237	=>	"000000000000000000000000000000",
1238	=>	"000000000000000000000000000000",
1239	=>	"000000000000000000000000000000",
1240	=>	"000000000000000000000000000000",
1241	=>	"000000000000000000000000000000",
1242	=>	"000000000000000000000000000000",
1243	=>	"000000000000000000000000000000",
1244	=>	"000000000000000000000000000000",
1245	=>	"000000000000000000000000000000",
1246	=>	"000000000000000000000000000000",
1247	=>	"000000000000000000000000000000",
1248	=>	"000000000000000000000000000000",
1249	=>	"000000000000000000000000000000",
1250	=>	"000000000000000000000000000000",
1251	=>	"000000000000000000000000000000",
1252	=>	"000000000000000000000000000000",
1253	=>	"000000000000000000000000000000",
1254	=>	"000000000000000000000000000000",
1255	=>	"000000000000000000000000000000",
1256	=>	"000000000000000000000000000000",
1257	=>	"000000000000000000000000000000",
1258	=>	"000000000000000000000000000000",
1259	=>	"000000000000000000000000000000",
1260	=>	"000000000000000000000000000000",
1261	=>	"000000000000000000000000000000",
1262	=>	"000000000000000000000000000000",
1263	=>	"000000000000000000000000000000",
1264	=>	"000000000000000000000000000000",
1265	=>	"000000000000000000000000000000",
1266	=>	"000000000000000000000000000000",
1267	=>	"000000000000000000000000000000",
1268	=>	"000000000000000000000000000000",
1269	=>	"000000000000000000000000000000",
1270	=>	"000000000000000000000000000000",
1271	=>	"000000000000000000000000000000",
1272	=>	"000000000000000000000000000000",
1273	=>	"000000000000000000000000000000",
1274	=>	"000000000000000000000000000000",
1275	=>	"000000000000000000000000000000",
1276	=>	"000000000000000000000000000000",
1277	=>	"000000000000000000000000000000",
1278	=>	"000000000000000000000000000000",
1279	=>	"000000000000000000000000000000",
1280	=>	"000000000000000000000000000000",
1281	=>	"000000000000000000000000000000",
1282	=>	"000000000000000000000000000000",
1283	=>	"000000000000000000000000000000",
1284	=>	"000000000000000000000000000000",
1285	=>	"000000000000000000000000000000",
1286	=>	"000000000000000000000000000000",
1287	=>	"000000000000000000000000000000",
1288	=>	"000000000000000000000000000000",
1289	=>	"000000000000000000000000000000",
1290	=>	"000000000000000000000000000000",
1291	=>	"000000000000000000000000000000",
1292	=>	"000000000000000000000000000000",
1293	=>	"000000000000000000000000000000",
1294	=>	"000000000000000000000000000000",
1295	=>	"000000000000000000000000000000",
1296	=>	"000000000000000000000000000000",
1297	=>	"000000000000000000000000000000",
1298	=>	"000000000000000000000000000000",
1299	=>	"000000000000000000000000000000",
1300	=>	"000000000000000000000000000000",
1301	=>	"000000000000000000000000000000",
1302	=>	"000000000000000000000000000000",
1303	=>	"000000000000000000000000000000",
1304	=>	"000000000000000000000000000000",
1305	=>	"000000000000000000000000000000",
1306	=>	"000000000000000000000000000000",
1307	=>	"000000000000000000000000000000",
1308	=>	"000000000000000000000000000000",
1309	=>	"000000000000000000000000000000",
1310	=>	"000000000000000000000000000000",
1311	=>	"000000000000000000000000000000",
1312	=>	"000000000000000000000000000000",
1313	=>	"000000000000000000000000000000",
1314	=>	"000000000000000000000000000000",
1315	=>	"000000000000000000000000000000",
1316	=>	"000000000000000000000000000000",
1317	=>	"000000000000000000000000000000",
1318	=>	"000000000000000000000000000000",
1319	=>	"000000000000000000000000000000",
1320	=>	"000000000000000000000000000000",
1321	=>	"000000000000000000000000000000",
1322	=>	"000000000000000000000000000000",
1323	=>	"000000000000000000000000000000",
1324	=>	"000000000000000000000000000000",
1325	=>	"000000000000000000000000000000",
1326	=>	"000000000000000000000000000000",
1327	=>	"000000000000000000000000000000",
1328	=>	"000000000000000000000000000000",
1329	=>	"000000000000000000000000000000",
1330	=>	"000000000000000000000000000000",
1331	=>	"000000000000000000000000000000",
1332	=>	"000000000000000000000000000000",
1333	=>	"000000000000000000000000000000",
1334	=>	"000000000000000000000000000000",
1335	=>	"000000000000000000000000000000",
1336	=>	"000000000000000000000000000000",
1337	=>	"000000000000000000000000000000",
1338	=>	"000000000000000000000000000000",
1339	=>	"000000000000000000000000000000",
1340	=>	"000000000000000000000000000000",
1341	=>	"000000000000000000000000000000",
1342	=>	"000000000000000000000000000000",
1343	=>	"000000000000000000000000000000",
1344	=>	"000000000000000000000000000000",
1345	=>	"000000000000000000000000000000",
1346	=>	"000000000000000000000000000000",
1347	=>	"000000000000000000000000000000",
1348	=>	"000000000000000000000000000000",
1349	=>	"000000000000000000000000000000",
1350	=>	"000000000000000000000000000000",
1351	=>	"000000000000000000000000000000",
1352	=>	"000000000000000000000000000000",
1353	=>	"000000000000000000000000000000",
1354	=>	"000000000000000000000000000000",
1355	=>	"000000000000000000000000000000",
1356	=>	"000000000000000000000000000000",
1357	=>	"000000000000000000000000000000",
1358	=>	"000000000000000000000000000000",
1359	=>	"000000000000000000000000000000",
1360	=>	"000000000000000000000000000000",
1361	=>	"000000000000000000000000000000",
1362	=>	"000000000000000000000000000000",
1363	=>	"000000000000000000000000000000",
1364	=>	"000000000000000000000000000000",
1365	=>	"000000000000000000000000000000",
1366	=>	"000000000000000000000000000000",
1367	=>	"000000000000000000000000000000",
1368	=>	"000000000000000000000000000000",
1369	=>	"000000000000000000000000000000",
1370	=>	"000000000000000000000000000000",
1371	=>	"000000000000000000000000000000",
1372	=>	"000000000000000000000000000000",
1373	=>	"000000000000000000000000000000",
1374	=>	"000000000000000000000000000000",
1375	=>	"000000000000000000000000000000",
1376	=>	"000000000000000000000000000000",
1377	=>	"000000000000000000000000000000",
1378	=>	"000000000000000000000000000000",
1379	=>	"000000000000000000000000000000",
1380	=>	"000000000000000000000000000000",
1381	=>	"000000000000000000000000000000",
1382	=>	"000000000000000000000000000000",
1383	=>	"000000000000000000000000000000",
1384	=>	"000000000000000000000000000000",
1385	=>	"000000000000000000000000000000",
1386	=>	"000000000000000000000000000000",
1387	=>	"000000000000000000000000000000",
1388	=>	"000000000000000000000000000000",
1389	=>	"000000000000000000000000000000",
1390	=>	"000000000000000000000000000000",
1391	=>	"000000000000000000000000000000",
1392	=>	"000000000000000000000000000000",
1393	=>	"000000000000000000000000000000",
1394	=>	"000000000000000000000000000000",
1395	=>	"000000000000000000000000000000",
1396	=>	"000000000000000000000000000000",
1397	=>	"000000000000000000000000000000",
1398	=>	"000000000000000000000000000000",
1399	=>	"000000000000000000000000000000",
1400	=>	"000000000000000000000000000000",
1401	=>	"000000000000000000000000000000",
1402	=>	"000000000000000000000000000000",
1403	=>	"000000000000000000000000000000",
1404	=>	"000000000000000000000000000000",
1405	=>	"000000000000000000000000000000",
1406	=>	"000000000000000000000000000000",
1407	=>	"000000000000000000000000000000",
1408	=>	"000000000000000000000000000000",
1409	=>	"000000000000000000000000000000",
1410	=>	"000000000000000000000000000000",
1411	=>	"000000000000000000000000000000",
1412	=>	"000000000000000000000000000000",
1413	=>	"000000000000000000000000000000",
1414	=>	"000000000000000000000000000000",
1415	=>	"000000000000000000000000000000",
1416	=>	"000000000000000000000000000000",
1417	=>	"000000000000000000000000000000",
1418	=>	"000000000000000000000000000000",
1419	=>	"000000000000000000000000000000",
1420	=>	"000000000000000000000000000000",
1421	=>	"000000000000000000000000000000",
1422	=>	"000000000000000000000000000000",
1423	=>	"000000000000000000000000000000",
1424	=>	"000000000000000000000000000000",
1425	=>	"000000000000000000000000000000",
1426	=>	"000000000000000000000000000000",
1427	=>	"000000000000000000000000000000",
1428	=>	"000000000000000000000000000000",
1429	=>	"000000000000000000000000000000",
1430	=>	"000000000000000000000000000000",
1431	=>	"000000000000000000000000000000",
1432	=>	"000000000000000000000000000000",
1433	=>	"000000000000000000000000000000",
1434	=>	"000000000000000000000000000000",
1435	=>	"000000000000000000000000000000",
1436	=>	"000000000000000000000000000000",
1437	=>	"000000000000000000000000000000",
1438	=>	"000000000000000000000000000000",
1439	=>	"000000000000000000000000000000",
1440	=>	"000000000000000000000000000000",
1441	=>	"000000000000000000000000000000",
1442	=>	"000000000000000000000000000000",
1443	=>	"000000000000000000000000000000",
1444	=>	"000000000000000000000000000000",
1445	=>	"000000000000000000000000000000",
1446	=>	"000000000000000000000000000000",
1447	=>	"000000000000000000000000000000",
1448	=>	"000000000000000000000000000000",
1449	=>	"000000000000000000000000000000",
1450	=>	"000000000000000000000000000000",
1451	=>	"000000000000000000000000000000",
1452	=>	"000000000000000000000000000000",
1453	=>	"000000000000000000000000000000",
1454	=>	"000000000000000000000000000000",
1455	=>	"000000000000000000000000000000",
1456	=>	"000000000000000000000000000000",
1457	=>	"000000000000000000000000000000",
1458	=>	"000000000000000000000000000000",
1459	=>	"000000000000000000000000000000",
1460	=>	"000000000000000000000000000000",
1461	=>	"000000000000000000000000000000",
1462	=>	"000000000000000000000000000000",
1463	=>	"000000000000000000000000000000",
1464	=>	"000000000000000000000000000000",
1465	=>	"000000000000000000000000000000",
1466	=>	"000000000000000000000000000000",
1467	=>	"000000000000000000000000000000",
1468	=>	"000000000000000000000000000000",
1469	=>	"000000000000000000000000000000",
1470	=>	"000000000000000000000000000000",
1471	=>	"000000000000000000000000000000",
1472	=>	"000000000000000000000000000000",
1473	=>	"000000000000000000000000000000",
1474	=>	"000000000000000000000000000000",
1475	=>	"000000000000000000000000000000",
1476	=>	"000000000000000000000000000000",
1477	=>	"000000000000000000000000000000",
1478	=>	"000000000000000000000000000000",
1479	=>	"000000000000000000000000000000",
1480	=>	"000000000000000000000000000000",
1481	=>	"000000000000000000000000000000",
1482	=>	"000000000000000000000000000000",
1483	=>	"000000000000000000000000000000",
1484	=>	"000000000000000000000000000000",
1485	=>	"000000000000000000000000000000",
1486	=>	"000000000000000000000000000000",
1487	=>	"000000000000000000000000000000",
1488	=>	"000000000000000000000000000000",
1489	=>	"000000000000000000000000000000",
1490	=>	"000000000000000000000000000000",
1491	=>	"000000000000000000000000000000",
1492	=>	"000000000000000000000000000000",
1493	=>	"000000000000000000000000000000",
1494	=>	"000000000000000000000000000000",
1495	=>	"000000000000000000000000000000",
1496	=>	"000000000000000000000000000000",
1497	=>	"000000000000000000000000000000",
1498	=>	"000000000000000000000000000000",
1499	=>	"000000000000000000000000000000",
1500	=>	"000000000000000000000000000000",
1501	=>	"000000000000000000000000000000",
1502	=>	"000000000000000000000000000000",
1503	=>	"000000000000000000000000000000",
1504	=>	"000000000000000000000000000000",
1505	=>	"000000000000000000000000000000",
1506	=>	"000000000000000000000000000000",
1507	=>	"000000000000000000000000000000",
1508	=>	"000000000000000000000000000000",
1509	=>	"000000000000000000000000000000",
1510	=>	"000000000000000000000000000000",
1511	=>	"000000000000000000000000000000",
1512	=>	"000000000000000000000000000000",
1513	=>	"000000000000000000000000000000",
1514	=>	"000000000000000000000000000000",
1515	=>	"000000000000000000000000000000",
1516	=>	"000000000000000000000000000000",
1517	=>	"000000000000000000000000000000",
1518	=>	"000000000000000000000000000000",
1519	=>	"000000000000000000000000000000",
1520	=>	"000000000000000000000000000000",
1521	=>	"000000000000000000000000000000",
1522	=>	"000000000000000000000000000000",
1523	=>	"000000000000000000000000000000",
1524	=>	"000000000000000000000000000000",
1525	=>	"000000000000000000000000000000",
1526	=>	"000000000000000000000000000000",
1527	=>	"000000000000000000000000000000",
1528	=>	"000000000000000000000000000000",
1529	=>	"000000000000000000000000000000",
1530	=>	"000000000000000000000000000000",
1531	=>	"000000000000000000000000000000",
1532	=>	"000000000000000000000000000000",
1533	=>	"000000000000000000000000000000",
1534	=>	"000000000000000000000000000000",
1535	=>	"000000000000000000000000000000",
1536	=>	"000000000000000000000000000000",
1537	=>	"000000000000000000000000000000",
1538	=>	"000000000000000000000000000000",
1539	=>	"000000000000000000000000000000",
1540	=>	"000000000000000000000000000000",
1541	=>	"000000000000000000000000000000",
1542	=>	"000000000000000000000000000000",
1543	=>	"000000000000000000000000000000",
1544	=>	"000000000000000000000000000000",
1545	=>	"000000000000000000000000000000",
1546	=>	"000000000000000000000000000000",
1547	=>	"000000000000000000000000000000",
1548	=>	"000000000000000000000000000000",
1549	=>	"000000000000000000000000000000",
1550	=>	"000000000000000000000000000000",
1551	=>	"000000000000000000000000000000",
1552	=>	"000000000000000000000000000000",
1553	=>	"000000000000000000000000000000",
1554	=>	"000000000000000000000000000000",
1555	=>	"000000000000000000000000000000",
1556	=>	"000000000000000000000000000000",
1557	=>	"000000000000000000000000000000",
1558	=>	"000000000000000000000000000000",
1559	=>	"000000000000000000000000000000",
1560	=>	"000000000000000000000000000000",
1561	=>	"000000000000000000000000000000",
1562	=>	"000000000000000000000000000000",
1563	=>	"000000000000000000000000000000",
1564	=>	"000000000000000000000000000000",
1565	=>	"000000000000000000000000000000",
1566	=>	"000000000000000000000000000000",
1567	=>	"000000000000000000000000000000",
1568	=>	"000000000000000000000000000000",
1569	=>	"000000000000000000000000000000",
1570	=>	"000000000000000000000000000000",
1571	=>	"000000000000000000000000000000",
1572	=>	"000000000000000000000000000000",
1573	=>	"000000000000000000000000000000",
1574	=>	"000000000000000000000000000000",
1575	=>	"000000000000000000000000000000",
1576	=>	"000000000000000000000000000000",
1577	=>	"000000000000000000000000000000",
1578	=>	"000000000000000000000000000000",
1579	=>	"000000000000000000000000000000",
1580	=>	"000000000000000000000000000000",
1581	=>	"000000000000000000000000000000",
1582	=>	"000000000000000000000000000000",
1583	=>	"000000000000000000000000000000",
1584	=>	"000000000000000000000000000000",
1585	=>	"000000000000000000000000000000",
1586	=>	"000000000000000000000000000000",
1587	=>	"000000000000000000000000000000",
1588	=>	"000000000000000000000000000000",
1589	=>	"000000000000000000000000000000",
1590	=>	"000000000000000000000000000000",
1591	=>	"000000000000000000000000000000",
1592	=>	"000000000000000000000000000000",
1593	=>	"000000000000000000000000000000",
1594	=>	"000000000000000000000000000000",
1595	=>	"000000000000000000000000000000",
1596	=>	"000000000000000000000000000000",
1597	=>	"000000000000000000000000000000",
1598	=>	"000000000000000000000000000000",
1599	=>	"000000000000000000000000000000",
1600	=>	"000000000000000000000000000000",
1601	=>	"000000000000000000000000000000",
1602	=>	"000000000000000000000000000000",
1603	=>	"000000000000000000000000000000",
1604	=>	"000000000000000000000000000000",
1605	=>	"000000000000000000000000000000",
1606	=>	"000000000000000000000000000000",
1607	=>	"000000000000000000000000000000",
1608	=>	"000000000000000000000000000000",
1609	=>	"000000000000000000000000000000",
1610	=>	"000000000000000000000000000000",
1611	=>	"000000000000000000000000000000",
1612	=>	"000000000000000000000000000000",
1613	=>	"000000000000000000000000000000",
1614	=>	"000000000000000000000000000000",
1615	=>	"000000000000000000000000000000",
1616	=>	"000000000000000000000000000000",
1617	=>	"000000000000000000000000000000",
1618	=>	"000000000000000000000000000000",
1619	=>	"000000000000000000000000000000",
1620	=>	"000000000000000000000000000000",
1621	=>	"000000000000000000000000000000",
1622	=>	"000000000000000000000000000000",
1623	=>	"000000000000000000000000000000",
1624	=>	"000000000000000000000000000000",
1625	=>	"000000000000000000000000000000",
1626	=>	"000000000000000000000000000000",
1627	=>	"000000000000000000000000000000",
1628	=>	"000000000000000000000000000000",
1629	=>	"000000000000000000000000000000",
1630	=>	"000000000000000000000000000000",
1631	=>	"000000000000000000000000000000",
1632	=>	"000000000000000000000000000000",
1633	=>	"000000000000000000000000000000",
1634	=>	"000000000000000000000000000000",
1635	=>	"000000000000000000000000000000",
1636	=>	"000000000000000000000000000000",
1637	=>	"000000000000000000000000000000",
1638	=>	"000000000000000000000000000000",
1639	=>	"000000000000000000000000000000",
1640	=>	"000000000000000000000000000000",
1641	=>	"000000000000000000000000000000",
1642	=>	"000000000000000000000000000000",
1643	=>	"000000000000000000000000000000",
1644	=>	"000000000000000000000000000000",
1645	=>	"000000000000000000000000000000",
1646	=>	"000000000000000000000000000000",
1647	=>	"000000000000000000000000000000",
1648	=>	"000000000000000000000000000000",
1649	=>	"000000000000000000000000000000",
1650	=>	"000000000000000000000000000000",
1651	=>	"000000000000000000000000000000",
1652	=>	"000000000000000000000000000000",
1653	=>	"000000000000000000000000000000",
1654	=>	"000000000000000000000000000000",
1655	=>	"000000000000000000000000000000",
1656	=>	"000000000000000000000000000000",
1657	=>	"000000000000000000000000000000",
1658	=>	"000000000000000000000000000000",
1659	=>	"000000000000000000000000000000",
1660	=>	"000000000000000000000000000000",
1661	=>	"000000000000000000000000000000",
1662	=>	"000000000000000000000000000000",
1663	=>	"000000000000000000000000000000",
1664	=>	"000000000000000000000000000000",
1665	=>	"000000000000000000000000000000",
1666	=>	"000000000000000000000000000000",
1667	=>	"000000000000000000000000000000",
1668	=>	"000000000000000000000000000000",
1669	=>	"000000000000000000000000000000",
1670	=>	"000000000000000000000000000000",
1671	=>	"000000000000000000000000000000",
1672	=>	"000000000000000000000000000000",
1673	=>	"000000000000000000000000000000",
1674	=>	"000000000000000000000000000000",
1675	=>	"000000000000000000000000000000",
1676	=>	"000000000000000000000000000000",
1677	=>	"000000000000000000000000000000",
1678	=>	"000000000000000000000000000000",
1679	=>	"000000000000000000000000000000",
1680	=>	"000000000000000000000000000000",
1681	=>	"000000000000000000000000000000",
1682	=>	"000000000000000000000000000000",
1683	=>	"000000000000000000000000000000",
1684	=>	"000000000000000000000000000000",
1685	=>	"000000000000000000000000000000",
1686	=>	"000000000000000000000000000000",
1687	=>	"000000000000000000000000000000",
1688	=>	"000000000000000000000000000000",
1689	=>	"000000000000000000000000000000",
1690	=>	"000000000000000000000000000000",
1691	=>	"000000000000000000000000000000",
1692	=>	"000000000000000000000000000000",
1693	=>	"000000000000000000000000000000",
1694	=>	"000000000000000000000000000000",
1695	=>	"000000000000000000000000000000",
1696	=>	"000000000000000000000000000000",
1697	=>	"000000000000000000000000000000",
1698	=>	"000000000000000000000000000000",
1699	=>	"000000000000000000000000000000",
1700	=>	"000000000000000000000000000000",
1701	=>	"000000000000000000000000000000",
1702	=>	"000000000000000000000000000000",
1703	=>	"000000000000000000000000000000",
1704	=>	"000000000000000000000000000000",
1705	=>	"000000000000000000000000000000",
1706	=>	"000000000000000000000000000000",
1707	=>	"000000000000000000000000000000",
1708	=>	"000000000000000000000000000000",
1709	=>	"000000000000000000000000000000",
1710	=>	"000000000000000000000000000000",
1711	=>	"000000000000000000000000000000",
1712	=>	"000000000000000000000000000000",
1713	=>	"000000000000000000000000000000",
1714	=>	"000000000000000000000000000000",
1715	=>	"000000000000000000000000000000",
1716	=>	"000000000000000000000000000000",
1717	=>	"000000000000000000000000000000",
1718	=>	"000000000000000000000000000000",
1719	=>	"000000000000000000000000000000",
1720	=>	"000000000000000000000000000000",
1721	=>	"000000000000000000000000000000",
1722	=>	"000000000000000000000000000000",
1723	=>	"000000000000000000000000000000",
1724	=>	"000000000000000000000000000000",
1725	=>	"000000000000000000000000000000",
1726	=>	"000000000000000000000000000000",
1727	=>	"000000000000000000000000000000",
1728	=>	"000000000000000000000000000000",
1729	=>	"000000000000000000000000000000",
1730	=>	"000000000000000000000000000000",
1731	=>	"000000000000000000000000000000",
1732	=>	"000000000000000000000000000000",
1733	=>	"000000000000000000000000000000",
1734	=>	"000000000000000000000000000000",
1735	=>	"000000000000000000000000000000",
1736	=>	"000000000000000000000000000000",
1737	=>	"000000000000000000000000000000",
1738	=>	"000000000000000000000000000000",
1739	=>	"000000000000000000000000000000",
1740	=>	"000000000000000000000000000000",
1741	=>	"000000000000000000000000000000",
1742	=>	"000000000000000000000000000000",
1743	=>	"000000000000000000000000000000",
1744	=>	"000000000000000000000000000000",
1745	=>	"000000000000000000000000000000",
1746	=>	"000000000000000000000000000000",
1747	=>	"000000000000000000000000000000",
1748	=>	"000000000000000000000000000000",
1749	=>	"000000000000000000000000000000",
1750	=>	"000000000000000000000000000000",
1751	=>	"000000000000000000000000000000",
1752	=>	"000000000000000000000000000000",
1753	=>	"000000000000000000000000000000",
1754	=>	"000000000000000000000000000000",
1755	=>	"000000000000000000000000000000",
1756	=>	"000000000000000000000000000000",
1757	=>	"000000000000000000000000000000",
1758	=>	"000000000000000000000000000000",
1759	=>	"000000000000000000000000000000",
1760	=>	"000000000000000000000000000000",
1761	=>	"000000000000000000000000000000",
1762	=>	"000000000000000000000000000000",
1763	=>	"000000000000000000000000000000",
1764	=>	"000000000000000000000000000000",
1765	=>	"000000000000000000000000000000",
1766	=>	"000000000000000000000000000000",
1767	=>	"000000000000000000000000000000",
1768	=>	"000000000000000000000000000000",
1769	=>	"000000000000000000000000000000",
1770	=>	"000000000000000000000000000000",
1771	=>	"000000000000000000000000000000",
1772	=>	"000000000000000000000000000000",
1773	=>	"000000000000000000000000000000",
1774	=>	"000000000000000000000000000000",
1775	=>	"000000000000000000000000000000",
1776	=>	"000000000000000000000000000000",
1777	=>	"000000000000000000000000000000",
1778	=>	"000000000000000000000000000000",
1779	=>	"000000000000000000000000000000",
1780	=>	"000000000000000000000000000000",
1781	=>	"000000000000000000000000000000",
1782	=>	"000000000000000000000000000000",
1783	=>	"000000000000000000000000000000",
1784	=>	"000000000000000000000000000000",
1785	=>	"000000000000000000000000000000",
1786	=>	"000000000000000000000000000000",
1787	=>	"000000000000000000000000000000",
1788	=>	"000000000000000000000000000000",
1789	=>	"000000000000000000000000000000",
1790	=>	"000000000000000000000000000000",
1791	=>	"000000000000000000000000000000",
1792	=>	"000000000000000000000000000000",
1793	=>	"000000000000000000000000000000",
1794	=>	"000000000000000000000000000000",
1795	=>	"000000000000000000000000000000",
1796	=>	"000000000000000000000000000000",
1797	=>	"000000000000000000000000000000",
1798	=>	"000000000000000000000000000000",
1799	=>	"000000000000000000000000000000",
1800	=>	"000000000000000000000000000000",
1801	=>	"000000000000000000000000000000",
1802	=>	"000000000000000000000000000000",
1803	=>	"000000000000000000000000000000",
1804	=>	"000000000000000000000000000000",
1805	=>	"000000000000000000000000000000",
1806	=>	"000000000000000000000000000000",
1807	=>	"000000000000000000000000000000",
1808	=>	"000000000000000000000000000000",
1809	=>	"000000000000000000000000000000",
1810	=>	"000000000000000000000000000000",
1811	=>	"000000000000000000000000000000",
1812	=>	"000000000000000000000000000000",
1813	=>	"000000000000000000000000000000",
1814	=>	"000000000000000000000000000000",
1815	=>	"000000000000000000000000000000",
1816	=>	"000000000000000000000000000000",
1817	=>	"000000000000000000000000000000",
1818	=>	"000000000000000000000000000000",
1819	=>	"000000000000000000000000000000",
1820	=>	"000000000000000000000000000000",
1821	=>	"000000000000000000000000000000",
1822	=>	"000000000000000000000000000000",
1823	=>	"000000000000000000000000000000",
1824	=>	"000000000000000000000000000000",
1825	=>	"000000000000000000000000000000",
1826	=>	"000000000000000000000000000000",
1827	=>	"000000000000000000000000000000",
1828	=>	"000000000000000000000000000000",
1829	=>	"000000000000000000000000000000",
1830	=>	"000000000000000000000000000000",
1831	=>	"000000000000000000000000000000",
1832	=>	"000000000000000000000000000000",
1833	=>	"000000000000000000000000000000",
1834	=>	"000000000000000000000000000000",
1835	=>	"000000000000000000000000000000",
1836	=>	"000000000000000000000000000000",
1837	=>	"000000000000000000000000000000",
1838	=>	"000000000000000000000000000000",
1839	=>	"000000000000000000000000000000",
1840	=>	"000000000000000000000000000000",
1841	=>	"000000000000000000000000000000",
1842	=>	"000000000000000000000000000000",
1843	=>	"000000000000000000000000000000",
1844	=>	"000000000000000000000000000000",
1845	=>	"000000000000000000000000000000",
1846	=>	"000000000000000000000000000000",
1847	=>	"000000000000000000000000000000",
1848	=>	"000000000000000000000000000000",
1849	=>	"000000000000000000000000000000",
1850	=>	"000000000000000000000000000000",
1851	=>	"000000000000000000000000000000",
1852	=>	"000000000000000000000000000000",
1853	=>	"000000000000000000000000000000",
1854	=>	"000000000000000000000000000000",
1855	=>	"000000000000000000000000000000",
1856	=>	"000000000000000000000000000000",
1857	=>	"000000000000000000000000000000",
1858	=>	"000000000000000000000000000000",
1859	=>	"000000000000000000000000000000",
1860	=>	"000000000000000000000000000000",
1861	=>	"000000000000000000000000000000",
1862	=>	"000000000000000000000000000000",
1863	=>	"000000000000000000000000000000",
1864	=>	"000000000000000000000000000000",
1865	=>	"000000000000000000000000000000",
1866	=>	"000000000000000000000000000000",
1867	=>	"000000000000000000000000000000",
1868	=>	"000000000000000000000000000000",
1869	=>	"000000000000000000000000000000",
1870	=>	"000000000000000000000000000000",
1871	=>	"000000000000000000000000000000",
1872	=>	"000000000000000000000000000000",
1873	=>	"000000000000000000000000000000",
1874	=>	"000000000000000000000000000000",
1875	=>	"000000000000000000000000000000",
1876	=>	"000000000000000000000000000000",
1877	=>	"000000000000000000000000000000",
1878	=>	"000000000000000000000000000000",
1879	=>	"000000000000000000000000000000",
1880	=>	"000000000000000000000000000000",
1881	=>	"000000000000000000000000000000",
1882	=>	"000000000000000000000000000000",
1883	=>	"000000000000000000000000000000",
1884	=>	"000000000000000000000000000000",
1885	=>	"000000000000000000000000000000",
1886	=>	"000000000000000000000000000000",
1887	=>	"000000000000000000000000000000",
1888	=>	"000000000000000000000000000000",
1889	=>	"000000000000000000000000000000",
1890	=>	"000000000000000000000000000000",
1891	=>	"000000000000000000000000000000",
1892	=>	"000000000000000000000000000000",
1893	=>	"000000000000000000000000000000",
1894	=>	"000000000000000000000000000000",
1895	=>	"000000000000000000000000000000",
1896	=>	"000000000000000000000000000000",
1897	=>	"000000000000000000000000000000",
1898	=>	"000000000000000000000000000000",
1899	=>	"000000000000000000000000000000",
1900	=>	"000000000000000000000000000000",
1901	=>	"000000000000000000000000000000",
1902	=>	"000000000000000000000000000000",
1903	=>	"000000000000000000000000000000",
1904	=>	"000000000000000000000000000000",
1905	=>	"000000000000000000000000000000",
1906	=>	"000000000000000000000000000000",
1907	=>	"000000000000000000000000000000",
1908	=>	"000000000000000000000000000000",
1909	=>	"000000000000000000000000000000",
1910	=>	"000000000000000000000000000000",
1911	=>	"000000000000000000000000000000",
1912	=>	"000000000000000000000000000000",
1913	=>	"000000000000000000000000000000",
1914	=>	"000000000000000000000000000000",
1915	=>	"000000000000000000000000000000",
1916	=>	"000000000000000000000000000000",
1917	=>	"000000000000000000000000000000",
1918	=>	"000000000000000000000000000000",
1919	=>	"000000000000000000000000000000",
1920	=>	"000000000000000000000000000000",
1921	=>	"000000000000000000000000000000",
1922	=>	"000000000000000000000000000000",
1923	=>	"000000000000000000000000000000",
1924	=>	"000000000000000000000000000000",
1925	=>	"000000000000000000000000000000",
1926	=>	"000000000000000000000000000000",
1927	=>	"000000000000000000000000000000",
1928	=>	"000000000000000000000000000000",
1929	=>	"000000000000000000000000000000",
1930	=>	"000000000000000000000000000000",
1931	=>	"000000000000000000000000000000",
1932	=>	"000000000000000000000000000000",
1933	=>	"000000000000000000000000000000",
1934	=>	"000000000000000000000000000000",
1935	=>	"000000000000000000000000000000",
1936	=>	"000000000000000000000000000000",
1937	=>	"000000000000000000000000000000",
1938	=>	"000000000000000000000000000000",
1939	=>	"000000000000000000000000000000",
1940	=>	"000000000000000000000000000000",
1941	=>	"000000000000000000000000000000",
1942	=>	"000000000000000000000000000000",
1943	=>	"000000000000000000000000000000",
1944	=>	"000000000000000000000000000000",
1945	=>	"000000000000000000000000000000",
1946	=>	"000000000000000000000000000000",
1947	=>	"000000000000000000000000000000",
1948	=>	"000000000000000000000000000000",
1949	=>	"000000000000000000000000000000",
1950	=>	"000000000000000000000000000000",
1951	=>	"000000000000000000000000000000",
1952	=>	"000000000000000000000000000000",
1953	=>	"000000000000000000000000000000",
1954	=>	"000000000000000000000000000000",
1955	=>	"000000000000000000000000000000",
1956	=>	"000000000000000000000000000000",
1957	=>	"000000000000000000000000000000",
1958	=>	"000000000000000000000000000000",
1959	=>	"000000000000000000000000000000",
1960	=>	"000000000000000000000000000000",
1961	=>	"000000000000000000000000000000",
1962	=>	"000000000000000000000000000000",
1963	=>	"000000000000000000000000000000",
1964	=>	"000000000000000000000000000000",
1965	=>	"000000000000000000000000000000",
1966	=>	"000000000000000000000000000000",
1967	=>	"000000000000000000000000000000",
1968	=>	"000000000000000000000000000000",
1969	=>	"000000000000000000000000000000",
1970	=>	"000000000000000000000000000000",
1971	=>	"000000000000000000000000000000",
1972	=>	"000000000000000000000000000000",
1973	=>	"000000000000000000000000000000",
1974	=>	"000000000000000000000000000000",
1975	=>	"000000000000000000000000000000",
1976	=>	"000000000000000000000000000000",
1977	=>	"000000000000000000000000000000",
1978	=>	"000000000000000000000000000000",
1979	=>	"000000000000000000000000000000",
1980	=>	"000000000000000000000000000000",
1981	=>	"000000000000000000000000000000",
1982	=>	"000000000000000000000000000000",
1983	=>	"000000000000000000000000000000",
1984	=>	"000000000000000000000000000000",
1985	=>	"000000000000000000000000000000",
1986	=>	"000000000000000000000000000000",
1987	=>	"000000000000000000000000000000",
1988	=>	"000000000000000000000000000000",
1989	=>	"000000000000000000000000000000",
1990	=>	"000000000000000000000000000000",
1991	=>	"000000000000000000000000000000",
1992	=>	"000000000000000000000000000000",
1993	=>	"000000000000000000000000000000",
1994	=>	"000000000000000000000000000000",
1995	=>	"000000000000000000000000000000",
1996	=>	"000000000000000000000000000000",
1997	=>	"000000000000000000000000000000",
1998	=>	"000000000000000000000000000000",
1999	=>	"000000000000000000000000000000",
2000	=>	"000000000000000000000000000000",
2001	=>	"000000000000000000000000000000",
2002	=>	"000000000000000000000000000000",
2003	=>	"000000000000000000000000000000",
2004	=>	"000000000000000000000000000000",
2005	=>	"000000000000000000000000000000",
2006	=>	"000000000000000000000000000000",
2007	=>	"000000000000000000000000000000",
2008	=>	"000000000000000000000000000000",
2009	=>	"000000000000000000000000000000",
2010	=>	"000000000000000000000000000000",
2011	=>	"000000000000000000000000000000",
2012	=>	"000000000000000000000000000000",
2013	=>	"000000000000000000000000000000",
2014	=>	"000000000000000000000000000000",
2015	=>	"000000000000000000000000000000",
2016	=>	"000000000000000000000000000000",
2017	=>	"000000000000000000000000000000",
2018	=>	"000000000000000000000000000000",
2019	=>	"000000000000000000000000000000",
2020	=>	"000000000000000000000000000000",
2021	=>	"000000000000000000000000000000",
2022	=>	"000000000000000000000000000000",
2023	=>	"000000000000000000000000000000",
2024	=>	"000000000000000000000000000000",
2025	=>	"000000000000000000000000000000",
2026	=>	"000000000000000000000000000000",
2027	=>	"000000000000000000000000000000",
2028	=>	"000000000000000000000000000000",
2029	=>	"000000000000000000000000000000",
2030	=>	"000000000000000000000000000000",
2031	=>	"000000000000000000000000000000",
2032	=>	"000000000000000000000000000000",
2033	=>	"000000000000000000000000000000",
2034	=>	"000000000000000000000000000000",
2035	=>	"000000000000000000000000000000",
2036	=>	"000000000000000000000000000000",
2037	=>	"000000000000000000000000000000",
2038	=>	"000000000000000000000000000000",
2039	=>	"000000000000000000000000000000",
2040	=>	"000000000000000000000000000000",
2041	=>	"000000000000000000000000000000",
2042	=>	"000000000000000000000000000000",
2043	=>	"000000000000000000000000000000",
2044	=>	"000000000000000000000000000000",
2045	=>	"000000000000000000000000000000",
2046	=>	"000000000000000000000000000000",
2047	=>	"000000000000000000000000000000"
);


signal 	LUT_data : std_logic_vector(C_Size_ROM_Sig+C_Size_ROM_Delta-1 downto 0);
signal	Sig	: unsigned(C_Size_ROM_Sig-1 downto 0);
signal	Delta	: signed(C_Size_ROM_Delta-1 downto 0);
signal	Intrp : signed(C_Size_in-C_ROM_Depth-1+1 downto 0);	--+1 for the sign bit
signal	DeltIntrp : signed(Delta'length+Intrp'length-1 downto 0);
signal	Func_out_buf : signed(C_Size_out-1+1 downto 0);

begin

LUT_data <= cts_rom_data(to_integer(Func_in(C_Size_in-1 downto C_Size_in-C_ROM_Depth)));

Delta <= signed(LUT_data(C_Size_ROM_Delta-1 downto 0));
Intrp	<= signed('0' & Func_in(C_Size_in-C_ROM_Depth-1 downto 0));

P_readout: process (CLK,RESET)
begin
	if(RESET = '1') then
		Sig			<= (others=>'0');
		DeltIntrp	<= (others=>'0');
	elsif rising_edge(CLK) then
		if (ENABLE_CLK ='1') then
			Sig 		 <= unsigned(LUT_data(C_Size_ROM_Sig+C_Size_ROM_Delta-1 downto C_Size_ROM_Delta));
			DeltIntrp <= Delta*Intrp;
		end if;
	end if;
end process;

Func_out_buf 	<= resize(signed('0' & Sig) + DeltIntrp(DeltIntrp'length-2 downto DeltIntrp'length-C_Size_ROM_Delta-1),Func_out_buf'length);
Func_out		<= unsigned(Func_out_buf(Func_out_buf'length-2 downto 0));

end Behavioral;